<!DOCTYPE html>
<html lang="sv">
<head>
  <meta http-equiv="Content-Type" content="text/html;charset=utf-8" >
  <meta name="yandex-verification" content="52297d544556772d" />
  <meta name="google-site-verification" content="ah8fN8rvRWoqb1FzT4B-uAfR1MwRdWvYzhyAFKXFWS8" />
  <meta name="viewport" content="width=device-width, initial-scale=1">
  <!-- WT_021 -->
  <title>BallroomDJ 4 - Musikspelare för balsalar</title>
  <!-- WT_022 -->
  <meta name="Description" content="BallroomDJ 4 - Musikspelare för balsalar">
  <meta name="Keywords" content="Ballroom Music Player,
      Přehrávač taneční hudby,
      Ballroom musikafspiller,
      Ballroom-Musikspieler,
      Reproductor de música de salón,
      Ballroom-musiikkisoitin,
      Lecteur de musique de salon,
      Bálterem zene lejátszó,
      Lettore di musica da sala da ballo,
      ボールルーム・ミュージック・プレーヤー,
      볼룸 음악 플레이어,
      Ballroom Muziekspeler,
      Odtwarzacz muzyki z sali balowej,
      Leitor de música de salão,
      Ballroom Музыкальный плеер,
      Musikspelare för balsalar,
      програвач бальної музики,
      舞厅音乐播放器,
      舞廳音樂播放器,
      ballroom music dj, ballroom dance dj,
      ballroom music playback,
      ballroom dance software,
      ballroom dance music software,
      ballroom dj software, ballroom dance software,
      dance studio music software,
      dance school music software,
      tango music player, tango dance player,
      country music player, country dance player">
  <link rel="stylesheet" type="text/css" href="bdj4.css">
</head>
<body>
  <div class="dbgwhite">
    <div class="menuwidget">
      <!-- WT_023 -->
      <img src="/img/menu.svg"
          alt="Meny"
          onclick="javascript:setDisplay('menu');">
    </div>
    <div>
      <!-- WT_001 -->
      <img src="/img/ballroomdj4.svg"
        alt="BallroomDJ 4 - Musikspelaren för ballroom"
        width="50%" style="max-width: 420px">
    </div>
    <div class="donatewidget">
      <form action="https://www.paypal.com/cgi-bin/webscr" method="post" target="_blank">
        <input type="hidden" name="cmd" value="_s-xclick" />
        <input type="hidden" name="hosted_button_id" value="BLTFRDM5KHNDJ" />
        <input type="image" src="https://www.paypalobjects.com/en_US/i/btn/btn_donate_SM.gif" border="0" name="submit" title="PayPal - The safer, easier way to pay online!" alt="Donate with PayPal button" />
        <img alt="" border="0" src="https://www.paypal.com/en_US/i/scr/pixel.gif" width="1" height="1" />
      </form>
    </div>
  </div>
  <div>
    <div id="dmenu" class="mdiv dispnone divmenu">
      <div class="tleft dinlineblock">
        <ul id="" class="menu">
          <li id="" class="menuitem"
              onclick="javascript:setDisplay('bdj4');">BallroomDJ 4</li>
          <li id="" class="menuitem"
              onclick="javascript:setDisplay('bdj3');">BallroomDJ 3</li>
          <!-- WT_002 -->
          <li id="" class="menuitem"
              onclick="javascript:setDisplay('donate');">Donera</li>
        </ul>
      </div>
    </div>
    <div id="dbdj4" class="mdiv dispblock">
      <div class="dflex">
        <div class="tleft dtext">
          <!-- WT_003 -->
          <p>BallroomDJ 4 (BDJ4) är en musikspelare som är avsedd för stationära och bärbara datorer (och fungerar även på vissa surfplattor). Den är utformad för att kunna spela musik under hela kvällen utan att någon behöver ingripa.</p>
          <!-- WT_004 -->
          <p>BDJ4 är mycket anpassningsbart och ger möjlighet att organisera dansmusik och skapa låtlistor, automatiska spellistor och sekvenserade spellistor.</p>
          <!-- WT_005 -->
          <p>BDJ4 körs på Windows, MacOS och Linux.</p>
          <!-- WT_006 -->
          <p><b><a target="_blank"
              href="https://sourceforge.net/projects/ballroomdj4/files/"
              >Ladda ner BallroomDJ 4</a></b>&nbsp;&nbsp;&nbsp;(<span>senaste versionen</span> <b>#VERSION#</b>)</p>
          <!-- WT_007 -->
          <p><a target="_blank"
              href="https://sourceforge.net/p/ballroomdj4/wiki/en-Change%20Log"
              >Ändra logg</a></p>
          <!-- WT_008 -->
          <p><a target="_blank"
              href="https://ballroomdj.org/forum/">BDJ4 Forum</a></p>
          <!-- WT_009 -->
          <p><a target="_blank"
              href="https://sourceforge.net/p/ballroomdj4/wiki/Home/"
              >BDJ4 Wiki</a></p>
          <!-- WT_010 -->
          <p><a target="_blank"
              href="https://sourceforge.net/p/ballroomdj4/wiki/en-Features/"
              >BDJ4 Funktioner</a></p>
          <!-- WT_011 -->
          <p><a target="_blank"
              href="https://crowdin.com/project/ballroomdj-4"
              >Hjälp att översätta BallroomDJ 4</a></p>
          <!-- WT_012 -->
          <p>Andra webbplatser där BallroomDJ 4 utgivningsmeddelanden kan hittas:</p>
          <!-- WT_013 -->
          <p><a target="_blank"
              href="https://freshcode.club/projects/bdj4"
              >BDJ4 på freshcode.club</a></p>
          <!-- WT_014 -->
          <p><a target="_blank"
              href="https://www.pro-linux.de/cgi-bin/DBApp/check.cgi?ShowAppDetail.01.17981.100"
              >BallroomDJ på pro-linux.de</a>  (Deutsch)</p>
        </div>
        <div class="tleft dlang">
          <ul>
            <li><a href="index.html.cs">čeština</a></li>
            <li><a href="index.html.da">Dansk</a></li>
            <li><a href="index.html.de">Deutsch</a></li>
            <li><a href="index.html.en">English</a></li>
            <li><a href="index.html.es-ES">Español</a></li>
            <li><a href="index.html.fi">Suomi</a></li>
            <li><a href="index.html.fr">Français</a></li>
            <li><a href="index.html.hu">magyar</a></li>
            <li><a href="index.html.it">Italiano</a></li>
            <li><a href="index.html.ja">日本語</a></li>
            <li><a href="index.html.ko">한국어</a></li>
            <li><a href="index.html.nb-NO">norsk</a></li>
            <li><a href="index.html.nl">Nederlands</a></li>
            <li><a href="index.html.pl-PL">Polski</a></li>
            <li><a href="index.html.pt-PT">Português</a></li>
            <li><a href="index.html.ru">Русский</a></li>
            <li><a href="index.html.sv">Svenska</a></li>
            <li><a href="index.html.uk">Українська</a></li>
            <li><a href="index.html.zh-CN">简体中文</a></li>
            <li><a href="index.html.zh-TW">繁體中文</a></li>
          </ul>
        </div>
      </div>
    </div>

    <div id="dbdj3" class="mdiv dispnone">
      <div class="tleft dinlineblock">
        <!-- WT_015 -->
        <p>BallroomDJ var den tidigare musikspelaren för balsalar. Den stöds inte längre.</p>
        <!-- WT_016 -->
        <p>Alla användare av BallroomDJ uppmanas att konvertera till BallroomDJ 4</p>
        <!-- WT_017 -->
        <p><a target="_blank"
            href="https://sourceforge.net/projects/ballroomdj/files/"
            >Ladda ner BallroomDJ 3</a></p>
      </div>
    </div>

    <div id="ddonate" class="mdiv dispnone tleft">
      <!-- WT_018 -->
      <p>Donera till BDJ4</p>
      <form action="https://www.paypal.com/cgi-bin/webscr" method="post" target="_blank">
        <input type="hidden" name="cmd" value="_s-xclick" />
        <input type="hidden" name="hosted_button_id" value="BLTFRDM5KHNDJ" />
        <input type="image" src="https://www.paypalobjects.com/en_US/i/btn/btn_donate_SM.gif" border="0" name="submit" title="PayPal - The safer, easier way to pay online!" alt="Donate with PayPal button" />
        <img alt="" border="0" src="https://www.paypal.com/en_US/i/scr/pixel.gif" width="1" height="1" />
      </form>
      <!-- WT_019 -->
      <p>Donera till mjukvaruprojekt som BDJ4 använder:</p>
      <!-- WT_020 -->
      <p><a href="https://videolan.org">VLC</a> (donationsknappen längst upp)</p>
      <p><a href="https://curl.se/donation.html">Curl</a></p>
      <p><a href="https://www.msys2.org/#donations">MSYS2</a> (Windows)</p>
      <p><a href="https://ffmpeg.org/donations.html">ffmpeg</a></p>
    </div>
  </div>

  <script type="text/javascript">
//<![CDATA[
function setDisplay (id) {
  if (id != 'menu') {
    var dids = {menu:0, bdj4:0, bdj3:0, donate:0};
    for (var i in dids) {
      var o = document.getElementById ('d'+i);
      o.style.display = 'none';
    }
  }

  var o = document.getElementById ('d'+id);
  o.style.display = 'block';
}
//]]>
  </script>
</body>
</html>
